`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:51:04 04/08/2020
// Design Name:   v74x139
// Module Name:   /home/ise/ise_projects/v74x139/test.v
// Project Name:  v74x139
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: v74x139
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test;

	// Inputs
	reg G_L1;
	reg G_L2;
	reg A1;
	reg A2;
	reg B1;
	reg B2;

	// Outputs
	wire [3:0] Y_L1;
	wire [3:0] Y_L2;

	// Instantiate the Unit Under Test (UUT)
	v74x139 uut (
		.G_L1(G_L1), 
		.G_L2(G_L2), 
		.A1(A1), 
		.A2(A2), 
		.B1(B1), 
		.B2(B2), 
		.Y_L1(Y_L1), 
		.Y_L2(Y_L2)
	);

	initial begin
		// Initialize Inputs
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 0;

		// Wait 100 ns for global reset to finish

        
		// Add stimulus here
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 0;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 0;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 0;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 0;
		B1 = 1;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 0;
		B2 = 1;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 0;
		#20;
		G_L1 = 1;
		G_L2 = 1;
		A1 = 1;
		A2 = 1;
		B1 = 1;
		B2 = 1;
		#20;

	end
      
endmodule

