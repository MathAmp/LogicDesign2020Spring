`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   08:04:21 04/28/2020
// Design Name:   hw
// Module Name:   /home/ise/ise_projects/HW5/vtest.v
// Project Name:  HW5
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: hw
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module vtest;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	hw uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#50;
        
		// Add stimulus here
		

	end
      
endmodule

